library verilog;
use verilog.vl_types.all;
entity tb_traffic_controller_1 is
end tb_traffic_controller_1;
