library verilog;
use verilog.vl_types.all;
entity tb_traffic_controller is
end tb_traffic_controller;
